module MemoryStage(

);

    

endmodule